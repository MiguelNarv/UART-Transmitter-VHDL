LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY EvenParityGenerator IS 
	GENERIC(
	BUSWIDTH: integer:=8
	);
	PORT(
	DATA: IN std_logic_vector(BUSWIDTH-1 DOWNTO 0);
	PARITY: OUT std_logic
	);
END ENTITY EvenParityGenerator;


ARCHITECTURE DataFlow OF EvenParityGenerator IS

BEGIN
	
	WITH BUSWIDTH SELECT 
	PARITY<=(((DATA(0) XOR DATA(1))XOR(DATA(2) XOR DATA(3))) XOR ((DATA(4) XOR DATA(5))XOR(DATA(6) XOR DATA(7)))) WHEN 8,
			(((DATA(0) XOR DATA(1))XOR(DATA(2) XOR DATA(3))) XOR ((DATA(4) XOR DATA(5))XOR(DATA(6) XOR '0'))) WHEN OTHERS;
	
END ARCHITECTURE DataFlow;